`timescale 1ns/1ns
module d_ff (
    input clk,
    input d,
    input rst,
    output reg q,
    output reg qb
);
    always @(negedge clk or negedge rst) begin
        if (rst == 1'b0) begin
            q <= 1'b0;
            qb <= 1'b1;
        end
        else begin
            q <= d;
            qb <= ~d;
        end
    end

endmodule: d_ff
